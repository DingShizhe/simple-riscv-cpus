
//Content of section .text

mem[0] = 32'h00000013;	// 0x0
mem[1] = 32'h0080006f;	// 0x4
mem[2] = 32'hffffffff;	// 0x8
mem[3] = 32'h00001137;	// 0xc
mem[4] = 32'h80010113;	// 0x10
mem[5] = 32'h0a4000ef;	// 0x14
mem[6] = 32'h00002423;	// 0x18
mem[7] = 32'h0000006f;	// 0x1c
mem[8] = 32'hfd010113;	// 0x20
mem[9] = 32'h02812623;	// 0x24
mem[10] = 32'h03010413;	// 0x28
mem[11] = 32'hfca42e23;	// 0x2c
mem[12] = 32'hfdc42703;	// 0x30
mem[13] = 32'h00c00793;	// 0x34
mem[14] = 32'h06e7e063;	// 0x38
mem[15] = 32'hfdc42783;	// 0x3c
mem[16] = 32'h00279713;	// 0x40
mem[17] = 32'h15c00793;	// 0x44
mem[18] = 32'h00f707b3;	// 0x48
mem[19] = 32'h0007a783;	// 0x4c
mem[20] = 32'h00078067;	// 0x50
mem[21] = 32'hfe042623;	// 0x54
mem[22] = 32'h04c0006f;	// 0x58
mem[23] = 32'h00200793;	// 0x5c
mem[24] = 32'hfef42623;	// 0x60
mem[25] = 32'h0400006f;	// 0x64
mem[26] = 32'h00500793;	// 0x68
mem[27] = 32'hfef42623;	// 0x6c
mem[28] = 32'h0340006f;	// 0x70
mem[29] = 32'h00800793;	// 0x74
mem[30] = 32'hfef42623;	// 0x78
mem[31] = 32'h0280006f;	// 0x7c
mem[32] = 32'h00a00793;	// 0x80
mem[33] = 32'hfef42623;	// 0x84
mem[34] = 32'h01c0006f;	// 0x88
mem[35] = 32'h00f00793;	// 0x8c
mem[36] = 32'hfef42623;	// 0x90
mem[37] = 32'h0100006f;	// 0x94
mem[38] = 32'hfff00793;	// 0x98
mem[39] = 32'hfef42623;	// 0x9c
mem[40] = 32'h00000013;	// 0xa0
mem[41] = 32'hfec42783;	// 0xa4
mem[42] = 32'h00078513;	// 0xa8
mem[43] = 32'h02c12403;	// 0xac
mem[44] = 32'h03010113;	// 0xb0
mem[45] = 32'h00008067;	// 0xb4
mem[46] = 32'hfe010113;	// 0xb8
mem[47] = 32'h00112e23;	// 0xbc
mem[48] = 32'h00812c23;	// 0xc0
mem[49] = 32'h02010413;	// 0xc4
mem[50] = 32'hfe042623;	// 0xc8
mem[51] = 32'h0500006f;	// 0xcc
mem[52] = 32'hfec42783;	// 0xd0
mem[53] = 32'hfff78793;	// 0xd4
mem[54] = 32'h00078513;	// 0xd8
mem[55] = 32'hf45ff0ef;	// 0xdc
mem[56] = 32'h00050693;	// 0xe0
mem[57] = 32'h000017b7;	// 0xe4
mem[58] = 32'hfec42703;	// 0xe8
mem[59] = 32'h00271713;	// 0xec
mem[60] = 32'h19078793;	// 0xf0
mem[61] = 32'h00f707b3;	// 0xf4
mem[62] = 32'h0007a783;	// 0xf8
mem[63] = 32'h00f68a63;	// 0xfc
mem[64] = 32'h000007b7;	// 0x100
mem[65] = 32'h00100713;	// 0x104
mem[66] = 32'h00e7a423;	// 0x108
mem[67] = 32'hf11ff06f;	// 0x10c
mem[68] = 32'hfec42783;	// 0x110
mem[69] = 32'h00178793;	// 0x114
mem[70] = 32'hfef42623;	// 0x118
mem[71] = 32'hfec42703;	// 0x11c
mem[72] = 32'h00e00793;	// 0x120
mem[73] = 32'hfae7d6e3;	// 0x124
mem[74] = 32'hfec42703;	// 0x128
mem[75] = 32'h00f00793;	// 0x12c
mem[76] = 32'h00f70a63;	// 0x130
mem[77] = 32'h000007b7;	// 0x134
mem[78] = 32'h00100713;	// 0x138
mem[79] = 32'h00e7a423;	// 0x13c
mem[80] = 32'heddff06f;	// 0x140
mem[81] = 32'h00000793;	// 0x144
mem[82] = 32'h00078513;	// 0x148
mem[83] = 32'h01c12083;	// 0x14c
mem[84] = 32'h01812403;	// 0x150
mem[85] = 32'h02010113;	// 0x154
mem[86] = 32'h00008067;	// 0x158

//Content of section .data

mem[87] = 32'h00000054;	// 0x15c
mem[88] = 32'h0000005c;	// 0x160
mem[89] = 32'h00000068;	// 0x164
mem[90] = 32'h00000068;	// 0x168
mem[91] = 32'h00000074;	// 0x16c
mem[92] = 32'h00000074;	// 0x170
mem[93] = 32'h00000074;	// 0x174
mem[94] = 32'h00000074;	// 0x178
mem[95] = 32'h00000080;	// 0x17c
mem[96] = 32'h00000080;	// 0x180
mem[97] = 32'h00000080;	// 0x184
mem[98] = 32'h00000080;	// 0x188
mem[99] = 32'h0000008c;	// 0x18c

//Content of section .data

mem[100] = 32'hffffffff;	// 0x190
mem[101] = 32'h00000000;	// 0x194
mem[102] = 32'h00000002;	// 0x198
mem[103] = 32'h00000005;	// 0x19c
mem[104] = 32'h00000005;	// 0x1a0
mem[105] = 32'h00000008;	// 0x1a4
mem[106] = 32'h00000008;	// 0x1a8
mem[107] = 32'h00000008;	// 0x1ac
mem[108] = 32'h00000008;	// 0x1b0
mem[109] = 32'h0000000a;	// 0x1b4
mem[110] = 32'h0000000a;	// 0x1b8
mem[111] = 32'h0000000a;	// 0x1bc
mem[112] = 32'h0000000a;	// 0x1c0
mem[113] = 32'h0000000f;	// 0x1c4
mem[114] = 32'hffffffff;	// 0x1c8

//Content of section .comment

//....
