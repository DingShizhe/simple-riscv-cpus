
//Content of section .text

mem[0] = 32'h00000013;	// 0x0
mem[1] = 32'h0080006f;	// 0x4
mem[2] = 32'hffffffff;	// 0x8
mem[3] = 32'h00001137;	// 0xc
mem[4] = 32'h80010113;	// 0x10
mem[5] = 32'h00c000ef;	// 0x14
mem[6] = 32'h00002423;	// 0x18
mem[7] = 32'h0000006f;	// 0x1c
mem[8] = 32'hff010113;	// 0x20
mem[9] = 32'h00812623;	// 0x24
mem[10] = 32'h01010413;	// 0x28
mem[11] = 32'h000017b7;	// 0x2c
mem[12] = 32'h1a07a223;	// 0x30
mem[13] = 32'h000017b7;	// 0x34
mem[14] = 32'h1a478793;	// 0x38
mem[15] = 32'h00100713;	// 0x3c
mem[16] = 32'h00e7a223;	// 0x40
mem[17] = 32'h000017b7;	// 0x44
mem[18] = 32'h1a478793;	// 0x48
mem[19] = 32'h00200713;	// 0x4c
mem[20] = 32'h00e7a423;	// 0x50
mem[21] = 32'h000017b7;	// 0x54
mem[22] = 32'h1a478793;	// 0x58
mem[23] = 32'h00300713;	// 0x5c
mem[24] = 32'h00e7a623;	// 0x60
mem[25] = 32'h000017b7;	// 0x64
mem[26] = 32'h1a478793;	// 0x68
mem[27] = 32'h00400713;	// 0x6c
mem[28] = 32'h00e7a823;	// 0x70
mem[29] = 32'h000017b7;	// 0x74
mem[30] = 32'h1a478793;	// 0x78
mem[31] = 32'h00c7a703;	// 0x7c
mem[32] = 32'h000017b7;	// 0x80
mem[33] = 32'h1ae7a023;	// 0x84
mem[34] = 32'h000017b7;	// 0x88
mem[35] = 32'h1a07a703;	// 0x8c
mem[36] = 32'h000017b7;	// 0x90
mem[37] = 32'h1a478793;	// 0x94
mem[38] = 32'h00e7aa23;	// 0x98
mem[39] = 32'h000017b7;	// 0x9c
mem[40] = 32'h1a47a783;	// 0xa0
mem[41] = 32'h00078a63;	// 0xa4
mem[42] = 32'h000007b7;	// 0xa8
mem[43] = 32'h00100713;	// 0xac
mem[44] = 32'h00e7a423;	// 0xb0
mem[45] = 32'hf69ff06f;	// 0xb4
mem[46] = 32'h000017b7;	// 0xb8
mem[47] = 32'h1a478793;	// 0xbc
mem[48] = 32'h0047a703;	// 0xc0
mem[49] = 32'h00100793;	// 0xc4
mem[50] = 32'h00f70a63;	// 0xc8
mem[51] = 32'h000007b7;	// 0xcc
mem[52] = 32'h00100713;	// 0xd0
mem[53] = 32'h00e7a423;	// 0xd4
mem[54] = 32'hf45ff06f;	// 0xd8
mem[55] = 32'h000017b7;	// 0xdc
mem[56] = 32'h1a478793;	// 0xe0
mem[57] = 32'h0087a703;	// 0xe4
mem[58] = 32'h00200793;	// 0xe8
mem[59] = 32'h00f70a63;	// 0xec
mem[60] = 32'h000007b7;	// 0xf0
mem[61] = 32'h00100713;	// 0xf4
mem[62] = 32'h00e7a423;	// 0xf8
mem[63] = 32'hf21ff06f;	// 0xfc
mem[64] = 32'h000017b7;	// 0x100
mem[65] = 32'h1a478793;	// 0x104
mem[66] = 32'h00c7a703;	// 0x108
mem[67] = 32'h00300793;	// 0x10c
mem[68] = 32'h00f70a63;	// 0x110
mem[69] = 32'h000007b7;	// 0x114
mem[70] = 32'h00100713;	// 0x118
mem[71] = 32'h00e7a423;	// 0x11c
mem[72] = 32'hefdff06f;	// 0x120
mem[73] = 32'h000017b7;	// 0x124
mem[74] = 32'h1a478793;	// 0x128
mem[75] = 32'h0107a703;	// 0x12c
mem[76] = 32'h00400793;	// 0x130
mem[77] = 32'h00f70a63;	// 0x134
mem[78] = 32'h000007b7;	// 0x138
mem[79] = 32'h00100713;	// 0x13c
mem[80] = 32'h00e7a423;	// 0x140
mem[81] = 32'hed9ff06f;	// 0x144
mem[82] = 32'h000017b7;	// 0x148
mem[83] = 32'h1a07a703;	// 0x14c
mem[84] = 32'h00300793;	// 0x150
mem[85] = 32'h00f70a63;	// 0x154
mem[86] = 32'h000007b7;	// 0x158
mem[87] = 32'h00100713;	// 0x15c
mem[88] = 32'h00e7a423;	// 0x160
mem[89] = 32'heb9ff06f;	// 0x164
mem[90] = 32'h000017b7;	// 0x168
mem[91] = 32'h1a478793;	// 0x16c
mem[92] = 32'h0147a703;	// 0x170
mem[93] = 32'h00300793;	// 0x174
mem[94] = 32'h00f70a63;	// 0x178
mem[95] = 32'h000007b7;	// 0x17c
mem[96] = 32'h00100713;	// 0x180
mem[97] = 32'h00e7a423;	// 0x184
mem[98] = 32'he95ff06f;	// 0x188
mem[99] = 32'h00000793;	// 0x18c
mem[100] = 32'h00078513;	// 0x190
mem[101] = 32'h00c12403;	// 0x194
mem[102] = 32'h01010113;	// 0x198
mem[103] = 32'h00008067;	// 0x19c

//Content of section .comment

//....
