
//Content of section .text

mem[0] = 32'h00000013;	// 0x0
mem[1] = 32'h0080006f;	// 0x4
mem[2] = 32'hffffffff;	// 0x8
mem[3] = 32'h00001137;	// 0xc
mem[4] = 32'h80010113;	// 0x10
mem[5] = 32'h00c000ef;	// 0x14
mem[6] = 32'h00002423;	// 0x18
mem[7] = 32'h0000006f;	// 0x1c
mem[8] = 32'hfe010113;	// 0x20
mem[9] = 32'h00812e23;	// 0x24
mem[10] = 32'h02010413;	// 0x28
mem[11] = 32'h00200793;	// 0x2c
mem[12] = 32'hfef42623;	// 0x30
mem[13] = 32'h0a80006f;	// 0x34
mem[14] = 32'hfec42783;	// 0x38
mem[15] = 32'hfff78713;	// 0x3c
mem[16] = 32'h000017b7;	// 0x40
mem[17] = 32'h00271713;	// 0x44
mem[18] = 32'h11878793;	// 0x48
mem[19] = 32'h00f707b3;	// 0x4c
mem[20] = 32'h0007a703;	// 0x50
mem[21] = 32'hfec42783;	// 0x54
mem[22] = 32'hffe78693;	// 0x58
mem[23] = 32'h000017b7;	// 0x5c
mem[24] = 32'h00269693;	// 0x60
mem[25] = 32'h11878793;	// 0x64
mem[26] = 32'h00f687b3;	// 0x68
mem[27] = 32'h0007a783;	// 0x6c
mem[28] = 32'h00f70733;	// 0x70
mem[29] = 32'h000017b7;	// 0x74
mem[30] = 32'hfec42683;	// 0x78
mem[31] = 32'h00269693;	// 0x7c
mem[32] = 32'h11878793;	// 0x80
mem[33] = 32'h00f687b3;	// 0x84
mem[34] = 32'h00e7a023;	// 0x88
mem[35] = 32'h000017b7;	// 0x8c
mem[36] = 32'hfec42703;	// 0x90
mem[37] = 32'h00271713;	// 0x94
mem[38] = 32'h11878793;	// 0x98
mem[39] = 32'h00f707b3;	// 0x9c
mem[40] = 32'h0007a703;	// 0xa0
mem[41] = 32'h000017b7;	// 0xa4
mem[42] = 32'hfec42683;	// 0xa8
mem[43] = 32'h00269693;	// 0xac
mem[44] = 32'h1b878793;	// 0xb0
mem[45] = 32'h00f687b3;	// 0xb4
mem[46] = 32'h0007a783;	// 0xb8
mem[47] = 32'h00f70a63;	// 0xbc
mem[48] = 32'h000007b7;	// 0xc0
mem[49] = 32'h00100713;	// 0xc4
mem[50] = 32'h00e7a423;	// 0xc8
mem[51] = 32'hf51ff06f;	// 0xcc
mem[52] = 32'hfec42783;	// 0xd0
mem[53] = 32'h00178793;	// 0xd4
mem[54] = 32'hfef42623;	// 0xd8
mem[55] = 32'hfec42703;	// 0xdc
mem[56] = 32'h02700793;	// 0xe0
mem[57] = 32'hf4e7dae3;	// 0xe4
mem[58] = 32'hfec42703;	// 0xe8
mem[59] = 32'h02800793;	// 0xec
mem[60] = 32'h00f70a63;	// 0xf0
mem[61] = 32'h000007b7;	// 0xf4
mem[62] = 32'h00100713;	// 0xf8
mem[63] = 32'h00e7a423;	// 0xfc
mem[64] = 32'hf1dff06f;	// 0x100
mem[65] = 32'h00000793;	// 0x104
mem[66] = 32'h00078513;	// 0x108
mem[67] = 32'h01c12403;	// 0x10c
mem[68] = 32'h02010113;	// 0x110
mem[69] = 32'h00008067;	// 0x114

//Content of section .data

mem[70] = 32'h00000001;	// 0x118
mem[71] = 32'h00000001;	// 0x11c
mem[72] = 32'h00000000;	// 0x120
mem[73] = 32'h00000000;	// 0x124
mem[74] = 32'h00000000;	// 0x128
mem[75] = 32'h00000000;	// 0x12c
mem[76] = 32'h00000000;	// 0x130
mem[77] = 32'h00000000;	// 0x134
mem[78] = 32'h00000000;	// 0x138
mem[79] = 32'h00000000;	// 0x13c
mem[80] = 32'h00000000;	// 0x140
mem[81] = 32'h00000000;	// 0x144
mem[82] = 32'h00000000;	// 0x148
mem[83] = 32'h00000000;	// 0x14c
mem[84] = 32'h00000000;	// 0x150
mem[85] = 32'h00000000;	// 0x154
mem[86] = 32'h00000000;	// 0x158
mem[87] = 32'h00000000;	// 0x15c
mem[88] = 32'h00000000;	// 0x160
mem[89] = 32'h00000000;	// 0x164
mem[90] = 32'h00000000;	// 0x168
mem[91] = 32'h00000000;	// 0x16c
mem[92] = 32'h00000000;	// 0x170
mem[93] = 32'h00000000;	// 0x174
mem[94] = 32'h00000000;	// 0x178
mem[95] = 32'h00000000;	// 0x17c
mem[96] = 32'h00000000;	// 0x180
mem[97] = 32'h00000000;	// 0x184
mem[98] = 32'h00000000;	// 0x188
mem[99] = 32'h00000000;	// 0x18c
mem[100] = 32'h00000000;	// 0x190
mem[101] = 32'h00000000;	// 0x194
mem[102] = 32'h00000000;	// 0x198
mem[103] = 32'h00000000;	// 0x19c
mem[104] = 32'h00000000;	// 0x1a0
mem[105] = 32'h00000000;	// 0x1a4
mem[106] = 32'h00000000;	// 0x1a8
mem[107] = 32'h00000000;	// 0x1ac
mem[108] = 32'h00000000;	// 0x1b0
mem[109] = 32'h00000000;	// 0x1b4
mem[110] = 32'h00000001;	// 0x1b8
mem[111] = 32'h00000001;	// 0x1bc
mem[112] = 32'h00000002;	// 0x1c0
mem[113] = 32'h00000003;	// 0x1c4
mem[114] = 32'h00000005;	// 0x1c8
mem[115] = 32'h00000008;	// 0x1cc
mem[116] = 32'h0000000d;	// 0x1d0
mem[117] = 32'h00000015;	// 0x1d4
mem[118] = 32'h00000022;	// 0x1d8
mem[119] = 32'h00000037;	// 0x1dc
mem[120] = 32'h00000059;	// 0x1e0
mem[121] = 32'h00000090;	// 0x1e4
mem[122] = 32'h000000e9;	// 0x1e8
mem[123] = 32'h00000179;	// 0x1ec
mem[124] = 32'h00000262;	// 0x1f0
mem[125] = 32'h000003db;	// 0x1f4
mem[126] = 32'h0000063d;	// 0x1f8
mem[127] = 32'h00000a18;	// 0x1fc
mem[128] = 32'h00001055;	// 0x200
mem[129] = 32'h00001a6d;	// 0x204
mem[130] = 32'h00002ac2;	// 0x208
mem[131] = 32'h0000452f;	// 0x20c
mem[132] = 32'h00006ff1;	// 0x210
mem[133] = 32'h0000b520;	// 0x214
mem[134] = 32'h00012511;	// 0x218
mem[135] = 32'h0001da31;	// 0x21c
mem[136] = 32'h0002ff42;	// 0x220
mem[137] = 32'h0004d973;	// 0x224
mem[138] = 32'h0007d8b5;	// 0x228
mem[139] = 32'h000cb228;	// 0x22c
mem[140] = 32'h00148add;	// 0x230
mem[141] = 32'h00213d05;	// 0x234
mem[142] = 32'h0035c7e2;	// 0x238
mem[143] = 32'h005704e7;	// 0x23c
mem[144] = 32'h008cccc9;	// 0x240
mem[145] = 32'h00e3d1b0;	// 0x244
mem[146] = 32'h01709e79;	// 0x248
mem[147] = 32'h02547029;	// 0x24c
mem[148] = 32'h03c50ea2;	// 0x250
mem[149] = 32'h06197ecb;	// 0x254

//Content of section .comment

//....
