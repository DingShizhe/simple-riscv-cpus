
//Content of section .text

mem[0] = 32'h00000013;	// 0x0
mem[1] = 32'h0080006f;	// 0x4
mem[2] = 32'hffffffff;	// 0x8
mem[3] = 32'h00001137;	// 0xc
mem[4] = 32'h80010113;	// 0x10
mem[5] = 32'h00c000ef;	// 0x14
mem[6] = 32'h00002423;	// 0x18
mem[7] = 32'h0000006f;	// 0x1c
mem[8] = 32'hfe010113;	// 0x20
mem[9] = 32'h00812e23;	// 0x24
mem[10] = 32'h02010413;	// 0x28
mem[11] = 32'h00100793;	// 0x2c
mem[12] = 32'hfef42623;	// 0x30
mem[13] = 32'hfe042423;	// 0x34
mem[14] = 32'h0200006f;	// 0x38
mem[15] = 32'hfe842703;	// 0x3c
mem[16] = 32'hfec42783;	// 0x40
mem[17] = 32'h00f707b3;	// 0x44
mem[18] = 32'hfef42423;	// 0x48
mem[19] = 32'hfec42783;	// 0x4c
mem[20] = 32'h00178793;	// 0x50
mem[21] = 32'hfef42623;	// 0x54
mem[22] = 32'hfec42703;	// 0x58
mem[23] = 32'h06400793;	// 0x5c
mem[24] = 32'hfce7dee3;	// 0x60
mem[25] = 32'hfe842703;	// 0x64
mem[26] = 32'h000017b7;	// 0x68
mem[27] = 32'h3ba78793;	// 0x6c
mem[28] = 32'h00f70a63;	// 0x70
mem[29] = 32'h000007b7;	// 0x74
mem[30] = 32'h00100713;	// 0x78
mem[31] = 32'h00e7a423;	// 0x7c
mem[32] = 32'hf9dff06f;	// 0x80
mem[33] = 32'h00000793;	// 0x84
mem[34] = 32'h00078513;	// 0x88
mem[35] = 32'h01c12403;	// 0x8c
mem[36] = 32'h02010113;	// 0x90
mem[37] = 32'h00008067;	// 0x94

//Content of section .comment

//....
