
//Content of section .text

mem[0] = 32'h00000013;	// 0x0
mem[1] = 32'h0080006f;	// 0x4
mem[2] = 32'hffffffff;	// 0x8
mem[3] = 32'h00001137;	// 0xc
mem[4] = 32'h80010113;	// 0x10
mem[5] = 32'h054000ef;	// 0x14
mem[6] = 32'h00002423;	// 0x18
mem[7] = 32'h0000006f;	// 0x1c
mem[8] = 32'hfd010113;	// 0x20
mem[9] = 32'h02812623;	// 0x24
mem[10] = 32'h03010413;	// 0x28
mem[11] = 32'hfca42e23;	// 0x2c
mem[12] = 32'hfcb42c23;	// 0x30
mem[13] = 32'hfdc42703;	// 0x34
mem[14] = 32'hfd842783;	// 0x38
mem[15] = 32'h00e7d863;	// 0x3c
mem[16] = 32'hfdc42783;	// 0x40
mem[17] = 32'hfef42623;	// 0x44
mem[18] = 32'h00c0006f;	// 0x48
mem[19] = 32'hfd842783;	// 0x4c
mem[20] = 32'hfef42623;	// 0x50
mem[21] = 32'hfec42783;	// 0x54
mem[22] = 32'h00078513;	// 0x58
mem[23] = 32'h02c12403;	// 0x5c
mem[24] = 32'h03010113;	// 0x60
mem[25] = 32'h00008067;	// 0x64
mem[26] = 32'hfe010113;	// 0x68
mem[27] = 32'h00112e23;	// 0x6c
mem[28] = 32'h00812c23;	// 0x70
mem[29] = 32'h02010413;	// 0x74
mem[30] = 32'hfe042223;	// 0x78
mem[31] = 32'hfe042623;	// 0x7c
mem[32] = 32'h0c00006f;	// 0x80
mem[33] = 32'hfe042423;	// 0x84
mem[34] = 32'h0840006f;	// 0x88
mem[35] = 32'h000017b7;	// 0x8c
mem[36] = 32'hfec42703;	// 0x90
mem[37] = 32'h00271713;	// 0x94
mem[38] = 32'h18078793;	// 0x98
mem[39] = 32'h00f707b3;	// 0x9c
mem[40] = 32'h0007a683;	// 0xa0
mem[41] = 32'h000017b7;	// 0xa4
mem[42] = 32'hfe842703;	// 0xa8
mem[43] = 32'h00271713;	// 0xac
mem[44] = 32'h18078793;	// 0xb0
mem[45] = 32'h00f707b3;	// 0xb4
mem[46] = 32'h0007a783;	// 0xb8
mem[47] = 32'h00078593;	// 0xbc
mem[48] = 32'h00068513;	// 0xc0
mem[49] = 32'hf5dff0ef;	// 0xc4
mem[50] = 32'h00050613;	// 0xc8
mem[51] = 32'hfe442783;	// 0xcc
mem[52] = 32'h00178713;	// 0xd0
mem[53] = 32'hfee42223;	// 0xd4
mem[54] = 32'h000016b7;	// 0xd8
mem[55] = 32'h00279713;	// 0xdc
mem[56] = 32'h1a068793;	// 0xe0
mem[57] = 32'h00f707b3;	// 0xe4
mem[58] = 32'h0007a783;	// 0xe8
mem[59] = 32'h00f60a63;	// 0xec
mem[60] = 32'h000007b7;	// 0xf0
mem[61] = 32'h00100713;	// 0xf4
mem[62] = 32'h00e7a423;	// 0xf8
mem[63] = 32'hf21ff06f;	// 0xfc
mem[64] = 32'hfe842783;	// 0x100
mem[65] = 32'h00178793;	// 0x104
mem[66] = 32'hfef42423;	// 0x108
mem[67] = 32'hfe842703;	// 0x10c
mem[68] = 32'h00700793;	// 0x110
mem[69] = 32'hf6e7fce3;	// 0x114
mem[70] = 32'hfe842703;	// 0x118
mem[71] = 32'h00800793;	// 0x11c
mem[72] = 32'h00f70a63;	// 0x120
mem[73] = 32'h000007b7;	// 0x124
mem[74] = 32'h00100713;	// 0x128
mem[75] = 32'h00e7a423;	// 0x12c
mem[76] = 32'heedff06f;	// 0x130
mem[77] = 32'hfec42783;	// 0x134
mem[78] = 32'h00178793;	// 0x138
mem[79] = 32'hfef42623;	// 0x13c
mem[80] = 32'hfec42703;	// 0x140
mem[81] = 32'h00700793;	// 0x144
mem[82] = 32'hf2e7fee3;	// 0x148
mem[83] = 32'hfec42703;	// 0x14c
mem[84] = 32'h00800793;	// 0x150
mem[85] = 32'h00f70a63;	// 0x154
mem[86] = 32'h000007b7;	// 0x158
mem[87] = 32'h00100713;	// 0x15c
mem[88] = 32'h00e7a423;	// 0x160
mem[89] = 32'heb9ff06f;	// 0x164
mem[90] = 32'h00000793;	// 0x168
mem[91] = 32'h00078513;	// 0x16c
mem[92] = 32'h01c12083;	// 0x170
mem[93] = 32'h01812403;	// 0x174
mem[94] = 32'h02010113;	// 0x178
mem[95] = 32'h00008067;	// 0x17c

//Content of section .data

mem[96] = 32'h00000000;	// 0x180
mem[97] = 32'h00000001;	// 0x184
mem[98] = 32'h00000002;	// 0x188
mem[99] = 32'h7fffffff;	// 0x18c
mem[100] = 32'h80000000;	// 0x190
mem[101] = 32'h80000001;	// 0x194
mem[102] = 32'hfffffffe;	// 0x198
mem[103] = 32'hffffffff;	// 0x19c
mem[104] = 32'h00000000;	// 0x1a0
mem[105] = 32'h00000001;	// 0x1a4
mem[106] = 32'h00000002;	// 0x1a8
mem[107] = 32'h7fffffff;	// 0x1ac
mem[108] = 32'h00000000;	// 0x1b0
mem[109] = 32'h00000000;	// 0x1b4
mem[110] = 32'h00000000;	// 0x1b8
mem[111] = 32'h00000000;	// 0x1bc
mem[112] = 32'h00000001;	// 0x1c0
mem[113] = 32'h00000001;	// 0x1c4
mem[114] = 32'h00000002;	// 0x1c8
mem[115] = 32'h7fffffff;	// 0x1cc
mem[116] = 32'h00000001;	// 0x1d0
mem[117] = 32'h00000001;	// 0x1d4
mem[118] = 32'h00000001;	// 0x1d8
mem[119] = 32'h00000001;	// 0x1dc
mem[120] = 32'h00000002;	// 0x1e0
mem[121] = 32'h00000002;	// 0x1e4
mem[122] = 32'h00000002;	// 0x1e8
mem[123] = 32'h7fffffff;	// 0x1ec
mem[124] = 32'h00000002;	// 0x1f0
mem[125] = 32'h00000002;	// 0x1f4
mem[126] = 32'h00000002;	// 0x1f8
mem[127] = 32'h00000002;	// 0x1fc
mem[128] = 32'h7fffffff;	// 0x200
mem[129] = 32'h7fffffff;	// 0x204
mem[130] = 32'h7fffffff;	// 0x208
mem[131] = 32'h7fffffff;	// 0x20c
mem[132] = 32'h7fffffff;	// 0x210
mem[133] = 32'h7fffffff;	// 0x214
mem[134] = 32'h7fffffff;	// 0x218
mem[135] = 32'h7fffffff;	// 0x21c
mem[136] = 32'h00000000;	// 0x220
mem[137] = 32'h00000001;	// 0x224
mem[138] = 32'h00000002;	// 0x228
mem[139] = 32'h7fffffff;	// 0x22c
mem[140] = 32'h80000000;	// 0x230
mem[141] = 32'h80000001;	// 0x234
mem[142] = 32'hfffffffe;	// 0x238
mem[143] = 32'hffffffff;	// 0x23c
mem[144] = 32'h00000000;	// 0x240
mem[145] = 32'h00000001;	// 0x244
mem[146] = 32'h00000002;	// 0x248
mem[147] = 32'h7fffffff;	// 0x24c
mem[148] = 32'h80000001;	// 0x250
mem[149] = 32'h80000001;	// 0x254
mem[150] = 32'hfffffffe;	// 0x258
mem[151] = 32'hffffffff;	// 0x25c
mem[152] = 32'h00000000;	// 0x260
mem[153] = 32'h00000001;	// 0x264
mem[154] = 32'h00000002;	// 0x268
mem[155] = 32'h7fffffff;	// 0x26c
mem[156] = 32'hfffffffe;	// 0x270
mem[157] = 32'hfffffffe;	// 0x274
mem[158] = 32'hfffffffe;	// 0x278
mem[159] = 32'hffffffff;	// 0x27c
mem[160] = 32'h00000000;	// 0x280
mem[161] = 32'h00000001;	// 0x284
mem[162] = 32'h00000002;	// 0x288
mem[163] = 32'h7fffffff;	// 0x28c
mem[164] = 32'hffffffff;	// 0x290
mem[165] = 32'hffffffff;	// 0x294
mem[166] = 32'hffffffff;	// 0x298
mem[167] = 32'hffffffff;	// 0x29c

//Content of section .comment

//....
